// $Id: $
// File name:   abc.sv
// Created:     9/15/2017
// Author:      Rtvik Sriram Bharadwaj
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: ksns.
